library verilog;
use verilog.vl_types.all;
entity decodModified_vlg_vec_tst is
end decodModified_vlg_vec_tst;
