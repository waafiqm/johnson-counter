library verilog;
use verilog.vl_types.all;
entity johnscirc_vlg_vec_tst is
end johnscirc_vlg_vec_tst;
