library verilog;
use verilog.vl_types.all;
entity muxModified_vlg_vec_tst is
end muxModified_vlg_vec_tst;
